/////////////////////////////////////////////////////////////////////////////////////
// 覴��ĵ㶥����ȡģ�飨ROM�������������棩
// �޸����ݣ�
// 1. ����ROM��λ���ԣ�active-high����ʹ��.rst(~rstn_out)
// 2. ��ַ��һ�ļĴ�(rom_addr_reg)������ͬ��ROMʱ��
// 3. �Ż�ROM���������߼���ȷ������ɼ����
// 4. ����ROM�������˿ڣ�tan_rom_addr/data/reg��cos_rom_addr/data/reg��
// 5. �޸��˿������﷨���ź���һ���Լ���λ��ʼ������
/////////////////////////////////////////////////////////////////////////////////////
module defect#(
    parameter IMG_WIDTH       = 11'd640,   // ͼ����
    parameter IMG_HEIGHT      = 11'd480,   // ͼ��߶�
    parameter COORD_WID       = 11,        // ����λ��0~2047��
    parameter TAN_REG_WID     = 16,        // tanֵ����Ĵ���λ����64�����ã�
    parameter ANGLE_WID       = 7,         // �Ƕ�λ��ƥ��ROM rd_data[6:0]��
    parameter DELAY_CYCLES    = 1,         // �ӳ�������1��2���ӳ٣�
    parameter SLOPE_THRESHOLD = 1,         // ��б�ж���ֵ
    parameter Z_DELTA_X       = 300        // ��������άz��Ƕ�
)(
    input                       pixclk_in,
    input                       rstn_out,   // �͵�ƽ��λ��ROM��λ�ź�ȡ��ʹ�ã�
    input                       bin2_vs,
    input                       bin2_de,
    input                       bin2_data,
    input                       set_template_flag,

    // ����������������ꡢ�������ꡢ��Ч��
    output reg [COORD_WID-1:0]  defect_p1_x,
    output reg [COORD_WID-1:0]  defect_p1_y,
    output reg [COORD_WID-1:0]  defect_p2_x,
    output reg [COORD_WID-1:0]  defect_p2_y,
    output reg [COORD_WID-1:0]  defect_p3_x,
    output reg [COORD_WID-1:0]  defect_p3_y,
    output reg [COORD_WID-1:0]  defect_p4_x,
    output reg [COORD_WID-1:0]  defect_p4_y,
    output reg [COORD_WID-1:0]  center_position_x,
    output reg [COORD_WID-1:0]  center_position_y,
    output reg                  defect_valid,
    output reg [ANGLE_WID-1:0]  angle,
    output reg [ANGLE_WID-1:0]  z_angle,
    output reg                  is_minus,   // 1Ϊ����0Ϊ��
    output                      point_vs,
    output                      point_de,

    // -------------------------- ������ROM�������˿� --------------------------
    // tan ROM��angle_rom���ӿ�
    output wire [11:0]          tan_rom_addr,      // ROM��ַ�������
    output wire [ANGLE_WID-1:0] tan_rom_data,      // ROMԭʼ���ݣ�δ���棬�����
    output reg [ANGLE_WID-1:0]  tan_rom_data_reg,  // ROM�������ݣ������
    // cos ROM��z_angle_rom���ӿ�
    output wire [11:0]          cos_rom_addr,      // ROM��ַ�������
    output wire [ANGLE_WID-1:0] cos_rom_data,      // ROMԭʼ���ݣ�δ���棬�����
    output reg [ANGLE_WID-1:0]  cos_rom_data_reg   // ROM�������ݣ������
    // --------------------------------------------------------------------------
);


/////////////////////////////////////////////////////////////////////////////////////
// 1. ���м�������ͼ�����������
/////////////////////////////////////////////////////////////////////////////////////
reg [COORD_WID-1:0] x_cnt, y_cnt;
always@(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        x_cnt <= 0;
    else if(x_cnt == IMG_WIDTH - 1'b1)
        x_cnt <= 0;
    else if(bin2_de)
        x_cnt <= x_cnt + 1'b1;

always@(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        y_cnt <= 0;
    else if(y_cnt == IMG_HEIGHT - 1'b1 && x_cnt == IMG_WIDTH - 1'b1)
        y_cnt <= 0;
    else if(x_cnt == IMG_WIDTH - 1'b1)
        y_cnt <= y_cnt + 1'b1;

/////////////////////////////////////////////////////////////////////////////////////
// 2. ��ֵ����߼�����ȡȱ�ݵ�x/y��ֵ����Ӧ���꣩
/////////////////////////////////////////////////////////////////////////////////////
reg [COORD_WID-1:0] x_min_reg, x_min_y_min_reg, x_min_y_max_reg;
reg [COORD_WID-1:0] x_max_reg, x_max_y_min_reg, x_max_y_max_reg;
reg [COORD_WID-1:0] y_min_reg, y_min_x_min_reg, y_min_x_max_reg;
reg [COORD_WID-1:0] y_max_reg, y_max_x_min_reg, y_max_x_max_reg;

reg bin2_vs_prev;
wire bin2_vs_posedge = bin2_vs && !bin2_vs_prev;  // ��ͬ�������أ�֡��ʼ��
always@(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        bin2_vs_prev <= 0;
    else
        bin2_vs_prev <= bin2_vs;

always @(posedge pixclk_in or negedge rstn_out) begin
    if (!rstn_out) begin
        // ��λʱ��ʼ����ֵ��x_min�����x_max����С��ȷ����֡�ܸ��£�
        x_min_reg <= IMG_WIDTH - 1'b1;  x_min_y_min_reg <= IMG_HEIGHT - 1'b1;  x_min_y_max_reg <= 0;
        x_max_reg <= 0;                 x_max_y_min_reg <= IMG_HEIGHT - 1'b1;  x_max_y_max_reg <= 0;
        y_min_reg <= IMG_HEIGHT - 1'b1; y_min_x_min_reg <= IMG_WIDTH - 1'b1;   y_min_x_max_reg <= 0;
        y_max_reg <= 0;                 y_max_x_min_reg <= IMG_WIDTH - 1'b1;   y_max_x_max_reg <= 0;
    end 
    else if (bin2_vs_posedge) begin
        // ÿ֡��ʼ���ü�ֵ��׼����֡��⣩
        x_min_reg <= IMG_WIDTH - 1'b1;  x_min_y_min_reg <= IMG_HEIGHT - 1'b1;  x_min_y_max_reg <= 0;
        x_max_reg <= 0;                 x_max_y_min_reg <= IMG_HEIGHT - 1'b1;  x_max_y_max_reg <= 0;
        y_min_reg <= IMG_HEIGHT - 1'b1; y_min_x_min_reg <= IMG_WIDTH - 1'b1;   y_min_x_max_reg <= 0;
        y_max_reg <= 0;                 y_max_x_min_reg <= IMG_WIDTH - 1'b1;   y_max_x_max_reg <= 0;
    end 
    else if (bin2_de && bin2_data == 1'b1) begin
        // ��⵽ȱ�����أ�bin2_data=1��������x/y��ֵ����Ӧy/x����
        // ����x��Сֵ��x_min������Ӧy�ļ�ֵ
        if (x_cnt < x_min_reg) begin
            x_min_reg       <= x_cnt;
            x_min_y_min_reg <= y_cnt;
            x_min_y_max_reg <= y_cnt;
        end else if (x_cnt == x_min_reg) begin
            if (y_cnt < x_min_y_min_reg) x_min_y_min_reg <= y_cnt;
            if (y_cnt > x_min_y_max_reg) x_min_y_max_reg <= y_cnt;
        end

        // ����x���ֵ��x_max������Ӧy�ļ�ֵ
        if (x_cnt > x_max_reg) begin
            x_max_reg       <= x_cnt;
            x_max_y_min_reg <= y_cnt;
            x_max_y_max_reg <= y_cnt;
        end else if (x_cnt == x_max_reg) begin
            if (y_cnt < x_max_y_min_reg) x_max_y_min_reg <= y_cnt;
            if (y_cnt > x_max_y_max_reg) x_max_y_max_reg <= y_cnt;
        end

        // ����y��Сֵ��y_min������Ӧx�ļ�ֵ
        if (y_cnt < y_min_reg) begin
            y_min_reg       <= y_cnt;
            y_min_x_min_reg <= x_cnt;
            y_min_x_max_reg <= x_cnt;
        end else if (y_cnt == y_min_reg) begin
            if (x_cnt < y_min_x_min_reg) y_min_x_min_reg <= x_cnt;
            if (x_cnt > y_min_x_max_reg) y_min_x_max_reg <= x_cnt;
        end

        // ����y���ֵ��y_max������Ӧx�ļ�ֵ
        if (y_cnt > y_max_reg) begin
            y_max_reg       <= y_cnt;
            y_max_x_min_reg <= x_cnt;
            y_max_x_max_reg <= x_cnt;
        end else if (y_cnt == y_max_reg) begin
            if (x_cnt < y_max_x_min_reg) y_max_x_min_reg <= x_cnt;
            if (x_cnt > y_max_x_max_reg) y_max_x_max_reg <= x_cnt;
        end
    end
end

/////////////////////////////////////////////////////////////////////////////////////
// 3. �������� + tan/cosֵ���㣨ȱ����״�жϼ��ǶȲ������㣩
/////////////////////////////////////////////////////////////////////////////////////
wire frame_end_flag = (x_cnt == IMG_WIDTH - 1'b1) && (y_cnt == IMG_HEIGHT - 1'b1);  // ֡������־
wire frame_has_defect = (x_min_reg <= x_max_reg);  // ֡���Ƿ����ȱ�ݣ�x_min��x_max��

// ��Ե��б�жϣ�����ؼ���Ե�Ĳ�ֵ
wire [COORD_WID-1:0] y_min_edge_diff = (x_min_y_min_reg > x_max_y_min_reg) ? 
                                       (x_min_y_min_reg - x_max_y_min_reg) : 
                                       (x_max_y_min_reg - x_min_y_min_reg);
wire [COORD_WID-1:0] x_min_edge_diff = (y_min_x_min_reg > y_max_x_min_reg) ? 
                                       (y_min_x_min_reg - y_max_x_min_reg) : 
                                       (y_max_x_min_reg - y_min_x_min_reg);
wire [COORD_WID-1:0] x_max_edge_diff = (y_min_x_max_reg > y_max_x_max_reg) ? 
                                       (y_min_x_max_reg - y_max_x_max_reg) : 
                                       (y_max_x_max_reg - y_min_x_max_reg);

// ȱ����״���ֱࣨ��/�ڰ�/��͹��
wire is_stright = (y_min_edge_diff < SLOPE_THRESHOLD) && (x_min_edge_diff < SLOPE_THRESHOLD);  // ֱ��
wire is_in      = (x_min_reg <= 10) && (x_max_reg > 0);  // �ڰ���x_min������߽磩
wire is_out     = (x_max_reg >= 630) && (x_min_reg > 0); // ��͹��x_max�����ұ߽磩

// �ڲ��Ĵ������������ꡢ�������ꡢtan/cosֵ����Ч��
reg [COORD_WID-1:0] p1_x_reg, p1_y_reg, p2_x_reg, p2_y_reg;
reg [COORD_WID-1:0] p3_x_reg, p3_y_reg, p4_x_reg, p4_y_reg;
reg [COORD_WID-1:0] p_x_reg, p_y_reg;
reg [TAN_REG_WID-1:0] tan_thita_reg;   // tanֵ�Ĵ���������tan ROM��ַ��
reg [TAN_REG_WID-1:0] z_cos_thita_reg; // cosֵ�Ĵ���������cos ROM��ַ��
reg valid_reg;                         // ȱ����Ч�ԼĴ���
reg is_minus_reg;                      // ������־�Ĵ���

// ����x_min��y_min����ľ��뼰�����ֵ������tanֵ���㣩
wire signed [COORD_WID-1:0] dx_1 = x_min_reg - y_min_x_min_reg;
wire signed [COORD_WID-1:0] dy_1 = x_min_y_min_reg - y_min_reg;
wire [COORD_WID-1:0] abs_dx_1 = (dx_1 < 0) ? -dx_1 : dx_1;
wire [COORD_WID-1:0] abs_dy_1 = (dy_1 < 0) ? -dy_1 : dy_1;
wire [COORD_WID-1:0] max_v_1 = (abs_dx_1 > abs_dy_1) ? abs_dx_1 : abs_dy_1;
wire [COORD_WID-1:0] min_v_1 = (abs_dx_1 > abs_dy_1) ? abs_dy_1 : abs_dx_1;
wire [COORD_WID-1:0] distance_approx_1 = max_v_1 
                                       + (min_v_1 >> 2) 
                                       + (min_v_1 >> 3);

// ����x_max��y_min����ľ��뼰�����ֵ�����������жϣ�
wire signed [COORD_WID-1:0] dx_2 = x_max_reg - y_min_x_max_reg;
wire signed [COORD_WID-1:0] dy_2 = x_max_y_min_reg - y_min_reg;
wire [COORD_WID-1:0] abs_dx_2 = (dx_2 < 0) ? -dx_2 : dx_2;
wire [COORD_WID-1:0] abs_dy_2 = (dy_2 < 0) ? -dy_2 : dy_2;
wire [COORD_WID-1:0] max_v_2 = (abs_dx_2 > abs_dy_2) ? abs_dx_2 : abs_dy_2;
wire [COORD_WID-1:0] min_v_2 = (abs_dx_2 > abs_dy_2) ? abs_dy_2 : abs_dx_2;
wire [COORD_WID-1:0] distance_approx_2 = max_v_2 
                                       + (min_v_2 >> 2) 
                                       + (min_v_2 >> 3);

// tanֵ���㣨��64�Ŵ󣬱���С����ʧ��
wire [TAN_REG_WID-1:0] dy_mul_64 = (distance_approx_1 > distance_approx_2) ? (abs_dy_1 << 6) : (abs_dy_2 << 6);
wire [TAN_REG_WID-1:0] dx_mul     = (distance_approx_1 > distance_approx_2) ? abs_dx_1 : abs_dx_2;
wire is_minus_wire                = (distance_approx_1 > distance_approx_2) ? 1'b1 : 1'b0;  // ������־
wire [TAN_REG_WID-1:0] tan_thita  = (dx_mul == 0) ? 16'd4095 : (dy_mul_64 / dx_mul);  // dx=0ʱ�����������

// ���㵱ǰdelta_x�����ڵ�set_template_flag=1ʱ��Ϊ�³�����
wire [COORD_WID-1:0] delta_x_current = (distance_approx_1 > distance_approx_2) ? distance_approx_1 : distance_approx_2;

// -------------------------- ���������л��ĳ����Ĵ��� --------------------------
reg [COORD_WID-1:0] divisor_reg;  // �洢��ǰ������Ĭ��Z_DELTA_X���ɱ�delta_x_current���£�

// �����Ĵ��������߼���
// - set_template_flag=1������ǰdelta_x_current����divisor_reg�����³�����
// - set_template_flag=0�����ֳ������䣨Ĭ��Z_DELTA_X���ϴθ���ֵ��
always @(posedge pixclk_in or negedge rstn_out) begin
    if (!rstn_out) begin
        divisor_reg <= Z_DELTA_X;  // ��λʱ��ʼ��ΪĬ�ϳ���
    end else if (set_template_flag == 1'b1) begin
        divisor_reg <= delta_x_current;  // �����ź���Чʱ����������Ϊ��ǰdelta_x
    end
    // else�����ֲ��䣬��ʹ��Ĭ��ֵ���ϴθ��µ�ֵ
end

// cosֵ���㣨����ͶӰ���߳���

wire [20:0] delta_longside_mul_4096 = delta_x_current << 12;  // ��������Ϊ��ǰdelta_x����ֵ
wire [TAN_REG_WID-1:0] z_cos_thita = (divisor_reg == 0) ? 16'd0 : (delta_longside_mul_4096 / divisor_reg);

// ֡����ʱ���涥�����ꡢtan/cosֵ��ÿ֡����һ�Σ�
always @(posedge pixclk_in or negedge rstn_out) begin
    if (!rstn_out) begin
        // ��λ��ʼ�������ڲ��Ĵ��������ⲻ��̬��
        {p1_x_reg, p1_y_reg, p2_x_reg, p2_y_reg, p3_x_reg, p3_y_reg, p4_x_reg, p4_y_reg} <= 0;
        p_x_reg <= 0;  p_y_reg <= 0;  tan_thita_reg <= 0;  z_cos_thita_reg <= 0;
        valid_reg <= 0;  is_minus_reg <= 1'b1;
    end else if (frame_end_flag) begin
        // ֡����������ȱ����״���涥������
        if(is_stright)begin  // 
            p1_x_reg <= x_min_reg;        p1_y_reg <= x_min_y_min_reg;
            p2_x_reg <= x_max_reg;        p2_y_reg <= x_max_y_min_reg;
            p3_x_reg <= y_max_x_min_reg;  p3_y_reg <= y_max_reg;
            p4_x_reg <= y_max_x_max_reg;  p4_y_reg <= y_max_reg;
            is_minus_reg <= 1'b1;
            tan_thita_reg <= 16'd4095;    // ֱ��tanֵ�����
            z_cos_thita_reg <= z_cos_thita;
        end else if(is_in)begin  // 
            p1_x_reg <= x_min_reg;        p1_y_reg <= x_min_y_min_reg;
            p2_x_reg <= x_max_reg;        p2_y_reg <= x_max_y_min_reg;
            p3_x_reg <= x_min_reg;        p3_y_reg <= x_min_y_max_reg;
            p4_x_reg <= y_max_x_max_reg;  p4_y_reg <= y_max_reg;
            is_minus_reg <= 1'b1;
            tan_thita_reg <= 16'd0;       // �ڰ�tanֵ��0
            z_cos_thita_reg <= 16'd0;
        end else if(is_out)begin  // 
            p1_x_reg <= x_min_reg;        p1_y_reg <= x_min_y_min_reg;
            p2_x_reg <= x_max_reg;        p2_y_reg <= x_max_y_min_reg;
            p3_x_reg <= y_max_x_min_reg;  p3_y_reg <= y_max_reg;
            p4_x_reg <= x_max_reg;        p4_y_reg <= x_max_y_max_reg;
            is_minus_reg <= 1'b1;
            //tan_thita_reg <= tan_thita;    // ��������tanֵ
            //z_cos_thita_reg <= z_cos_thita;
        end else begin  // 
            p1_x_reg <= x_min_reg;        p1_y_reg <= x_min_y_min_reg;
            p2_x_reg <= x_max_reg;        p2_y_reg <= x_max_y_min_reg;
            p3_x_reg <= y_min_x_min_reg;  p3_y_reg <= y_min_reg;
            p4_x_reg <= y_max_x_max_reg;  p4_y_reg <= y_max_reg;
            is_minus_reg <= is_minus_wire; // ����������־
            tan_thita_reg <= tan_thita;    // ��������tanֵ
            z_cos_thita_reg <= z_cos_thita;
        end
        // ����ȱ���������꣨ȡx/y��ֵ���е㣩
        p_x_reg <= (x_max_reg + x_min_reg + 1) >> 1;
        p_y_reg <= (y_max_reg + y_min_reg + 1) >> 1;
        valid_reg <= frame_has_defect;  // ����ȱ����Ч��
    end
end

/////////////////////////////////////////////////////////////////////////////////////
// 4. tan ROM�ӿڣ�angle_rom������ַ���ɡ���������
/////////////////////////////////////////////////////////////////////////////////////
reg [11:0] rom_addr_reg;          // tan ROM��ַ�Ĵ�����12λ��ƥ��4096��ȣ�
wire [ANGLE_WID-1:0] rom_tan_data;// tan ROMԭʼ������ݣ�7λ����Ӧ0~89�㣩

// tan ROM��ַ���ɣ���tan_thita_regȡ��12λ������ROM��ȣ�
always @(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        rom_addr_reg <= 12'd0;
    else
        rom_addr_reg <= tan_thita_reg[11:0];

// ����tan ROM���Ϲ�ͬ��DRM Based ROM����������IP����һ�£�
angle_rom angle_rom_inst (
    .addr   (rom_addr_reg),    // ROM��ַ�����룩
    .clk    (pixclk_in),       // ʱ�ӣ���ģ��ʱ��ͬ����
    .rst    (~rstn_out),       // ROM��λ��active-high����ģ�鸴λ����ƥ�䣩
    .rd_data(rom_tan_data)     // ROM���������7λ�Ƕ�ֵ��
);

// tan ROM�������棨ͬ��ʱ�ӣ�ȷ�������ȶ���
always @(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        tan_rom_data_reg <= 7'd0;  // ��λʱ����������0
    else
        tan_rom_data_reg <= rom_tan_data;  // ÿʱ��������ROM���

/////////////////////////////////////////////////////////////////////////////////////
// 5. cos ROM�ӿڣ�z_angle_rom������ַ���ɡ���������
/////////////////////////////////////////////////////////////////////////////////////
reg [11:0] rom_addr_reg_zcos;     // cos ROM��ַ�Ĵ�����12λ��ƥ��4096��ȣ�
wire [ANGLE_WID-1:0] rom_cos_data;// cos ROMԭʼ������ݣ�7λ����Ӧ0~89�㣩

// cos ROM��ַ���ɣ���z_cos_thita_regȡ��12λ������ROM��ȣ�
always @(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        rom_addr_reg_zcos <= 12'd0;
    else
        rom_addr_reg_zcos <= z_cos_thita_reg[11:0];

// ����cos ROM���Ϲ�ͬ��DRM Based ROM����������IP����һ�£�
z_angle_rom z_angle_rom_inst (
    .addr   (rom_addr_reg_zcos),// ROM��ַ�����룩
    .clk    (pixclk_in),        // ʱ�ӣ���ģ��ʱ��ͬ����
    .rst    (~rstn_out),        // ROM��λ��active-high����ģ�鸴λ����ƥ�䣩
    .rd_data(rom_cos_data)      // ROM���������7λ�Ƕ�ֵ��
);

// cos ROM�������棨ͬ��ʱ�ӣ�ȷ�������ȶ���
always @(posedge pixclk_in or negedge rstn_out)
    if(!rstn_out)
        cos_rom_data_reg <= 7'd0;  // ��λʱ����������0
    else
        cos_rom_data_reg <= rom_cos_data;  // ÿʱ��������ROM���

/////////////////////////////////////////////////////////////////////////////////////
// 6. ROM����˿ڰ󶨣����ڲ��ź�ӳ�䵽ģ�������
/////////////////////////////////////////////////////////////////////////////////////
assign tan_rom_addr = rom_addr_reg;      // tan ROM��ַ �� ģ�����
assign tan_rom_data = rom_tan_data;      // tan ROMԭʼ���� �� ģ�����
assign cos_rom_addr = rom_addr_reg_zcos; // cos ROM��ַ �� ģ�����
assign cos_rom_data = rom_cos_data;      // cos ROMԭʼ���� �� ģ�����

/////////////////////////////////////////////////////////////////////////////////////
// 7. ���������ͬ�������ڲ��Ĵ���ֵӳ�䵽ģ�����������
/////////////////////////////////////////////////////////////////////////////////////
reg [DELAY_CYCLES:0] vs_delay_chain, de_delay_chain;  // ��/����ʹ���ӳ�����ͬ�������
always @(posedge pixclk_in or negedge rstn_out)
    if (!rstn_out) begin
        vs_delay_chain <= 0;
        de_delay_chain <= 0;
    end else begin
        // �ӳ�����ȷ�������ͼ��ʱ��ͬ�����ӳ�DELAY_CYCLES+1�ģ�
        vs_delay_chain <= {vs_delay_chain[DELAY_CYCLES-1:0], bin2_vs};
        de_delay_chain <= {de_delay_chain[DELAY_CYCLES-1:0], bin2_de};
    end

// ����������棨ÿʱ���ظ��£����ӳ���ʱ��ƥ�䣩
always @(posedge pixclk_in or negedge rstn_out)
    if (!rstn_out) begin
        // ��λʱ���������0
        {defect_p1_x, defect_p1_y, defect_p2_x, defect_p2_y,
         defect_p3_x, defect_p3_y, defect_p4_x, defect_p4_y} <= 0;
        center_position_x <= 0;  center_position_y <= 0;
        angle <= 0;  z_angle <= 0;  defect_valid <= 0;  is_minus <= 1'b1;
    end else begin
        // ӳ���ڲ�����Ķ��㡢��������
        {defect_p1_x, defect_p1_y} <= {p1_x_reg, p1_y_reg};
        {defect_p2_x, defect_p2_y} <= {p2_x_reg, p2_y_reg};
        {defect_p3_x, defect_p3_y} <= {p3_x_reg, p3_y_reg};
        {defect_p4_x, defect_p4_y} <= {p4_x_reg, p4_y_reg};
        center_position_x <= p_x_reg;
        center_position_y <= p_y_reg;
// �ؼ��޸ģ���ȱ�ݡ�ROM�Ƕȣ���ȱ�ݡ�ǿ��0��
        angle <= valid_reg ? tan_rom_data_reg : 7'd0;  // ��ȱ��ʱangle=0��
        z_angle <= valid_reg ? cos_rom_data_reg : 7'd0;  // ��ȱ��ʱz_angleҲ��0�㣨��ѡ��������
        // ӳ��ȱ����Ч�ԡ�������־
        defect_valid <= valid_reg;
        is_minus <= is_minus_reg; 
    end

// ͬ����ĳ�/����ʹ�����
assign point_vs = vs_delay_chain[DELAY_CYCLES];
assign point_de = de_delay_chain[DELAY_CYCLES];

endmodule