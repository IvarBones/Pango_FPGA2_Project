//��ֵ�˲�   delay 3clk
module median_filter_3x3(
    input wire           clk       ,
    input wire           rst_n     ,
    input wire           vsync_in  ,
    input wire           hsync_in  ,
    input wire           de_in     ,
   
    input wire    [7:0]  data11    , 
    input wire    [7:0]  data12    , 
    input wire    [7:0]  data13    ,
    input wire    [7:0]  data21    , 
    input wire    [7:0]  data22    , 
    input wire    [7:0]  data23    ,
    input wire    [7:0]  data31    , 
    input wire    [7:0]  data32    , 
    input wire    [7:0]  data33    ,
   
    output wire   [7:0]  target_data,
    output wire          vsync_out  ,
    output wire          hsync_out  ,
    output wire          de_out
);

//--------------------------------------------------------------------------------------
//FPGA Median Filter Sort order
//       Pixel -- Sort1 -- Sort2 -- Sort3
// [ P1  P2  P3 ]   [   Max1  Mid1   Min1 ]
// [ P4  P5  P6 ]   [   Max2  Mid2   Min2 ] [Max_min, Mid_mid, Min_max] mid_valid
// [ P7  P8  P9 ]   [   Max3  Mid3   Min3 ]

//reg define
reg [2:0]   vsync_in_r;
reg [2:0]   hsync_in_r;
reg [2:0]   de_in_r;
//wire define
wire [7:0] max_data1; 
wire [7:0] mid_data1; 
wire [7:0] min_data1;
wire [7:0] max_data2; 
wire [7:0] mid_data2; 
wire [7:0] min_data2;
wire [7:0] max_data3; 
wire [7:0] mid_data3; 
wire [7:0] min_data3;
wire [7:0] max_min_data; 
wire [7:0] mid_mid_data; 
wire [7:0] min_max_data;

//*****************************************************
//**                    main code
//*****************************************************

assign vsync_out = vsync_in_r[2];
assign hsync_out  = hsync_in_r[2];
assign de_out = de_in_r[2];

//Step1 ��stor3����������������
sort3  u_sort3_1(     //��һ����������
    .clk      (clk),
    .rst_n    (rst_n),
    
    .data1    (data11), 
    .data2    (data12), 
    .data3    (data13),
    
    .max_data (max_data1),
    .mid_data (mid_data1),
    .min_data (min_data1)
);

sort3  u_sort3_2(      //�ڶ�����������
    .clk      (clk),
    .rst_n    (rst_n),
        
    .data1    (data21), 
    .data2    (data22), 
    .data3    (data23),
    
    .max_data (max_data2),
    .mid_data (mid_data2),
    .min_data (min_data2)
);

sort3  u_sort3_3(      //��������������
    .clk      (clk),
    .rst_n    (rst_n),
        
    .data1    (data31), 
    .data2    (data32), 
    .data3    (data33),
    
    .max_data (max_data3),
    .mid_data (mid_data3),
    .min_data (min_data3)
);

//Step2 ����������ȡ�õ�������д���
sort3 u_sort3_4(        //ȡ�������ֵ����Сֵ
    .clk      (clk),
    .rst_n    (rst_n),
          
    .data1    (max_data1), 
    .data2    (max_data2), 
    .data3    (max_data3),
    
    .max_data (),
    .mid_data (),
    .min_data (max_min_data)
);

sort3 u_sort3_5(        //ȡ������ֵ����Сֵ
    .clk      (clk),
    .rst_n    (rst_n),
          
    .data1    (mid_data1), 
    .data2    (mid_data2), 
    .data3    (mid_data3),
    
    .max_data (),
    .mid_data (mid_mid_data),
    .min_data ()
);

sort3 u_sort3_6(        //ȡ������Сֵ�����ֵ
    .clk      (clk),
    .rst_n    (rst_n),
          
    .data1    (min_data1), 
    .data2    (min_data2), 
    .data3    (min_data3),
    
    .max_data (min_max_data),
    .mid_data (),
    .min_data ()
);

//step3 ��step2 �еõ�������ֵ���ٴ�ȡ��ֵ
sort3 u_sort3_7(
    .clk      (clk),
    .rst_n    (rst_n),
          
    .data1    (max_min_data), 
    .data2    (mid_mid_data), 
    .data3    (min_max_data),
    
    .max_data (),
    .mid_data (target_data),
    .min_data ()
);

//�ӳ��������ڽ���ͬ��
always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        vsync_in_r <= 0;
        hsync_in_r  <= 0;
        de_in_r <= 0;
    end
    else begin
        vsync_in_r <= {vsync_in_r[1:0],vsync_in};
        hsync_in_r  <= {hsync_in_r [1:0], hsync_in};
        de_in_r <= {de_in_r[1:0],de_in};
    end
end

endmodule 