// ��������ģ�飨�����̹�100Pro+���͵�ƽ��Ч��27MHzʱ�ӣ�20ms������
module key#(
    parameter DEBOUNCE_CNT = 20'd540000  // 27MHz * 20ms = 540000��������ֵ
)(
    input               sys_clk      ,  // ����ʱ�ӣ�27MHz�����Զ��㣩
    input               rst_in       ,  // ���븴λ���͵�ƽ��Ч�����Զ���rst_in��
    input               key_raw      ,  // ���룺ԭʼ�����źţ��͵�ƽ��Ч��
    output reg          key_press    ,  // ������������δ������ߵ�ƽ1��ʱ�����ڣ�
    output reg          key_state     // �����������ǰ״̬����=���£���=δ���£�
);

// 1. �����Ĵ���ͬ������������̬���������ź�ͬ����sys_clk��
reg key_sync1, key_sync2;
always @(posedge sys_clk or negedge rst_in) begin
    if (!rst_in) begin  // ��λʱ������Ĭ��δ���£�ͬ����Ϊ�ߵ�ƽ��
        key_sync1 <= 1'b1;
        key_sync2 <= 1'b1;
    end else begin
        key_sync1 <= key_raw;       // ��һ��ͬ��
        key_sync2 <= key_sync1;     // �ڶ���ͬ���������ȶ��İ����źţ�
    end
end

// 2. ��������������ⰴ���ȶ�״̬��
reg [19:0] debounce_cnt;  // 20λ�㹻�洢540000�����ֵ2^20=1,048,576��
always @(posedge sys_clk or negedge rst_in) begin
    if (!rst_in) begin
        debounce_cnt <= 20'd0;
    end else begin
        if (key_sync2 == 1'b1) begin  // ����δ���£��ߵ�ƽ��������������
            debounce_cnt <= 20'd0;
        end else begin  // �������£��͵�ƽ�����������ۼӣ�ֱ����ֵ
            debounce_cnt <= (debounce_cnt >= DEBOUNCE_CNT) ? DEBOUNCE_CNT : debounce_cnt + 1'b1;
        end
    end
end

// 3. ���ɰ���״̬�뵥�δ����ź�
reg debounce_cnt_prev;  // ��¼��һ���ڼ������Ƿ������������ɵ����ڴ���
always @(posedge sys_clk or negedge rst_in) begin
    if (!rst_in) begin
        key_state <= 1'b0;        // ��λʱ����δ����
        debounce_cnt_prev <= 1'b0;
        key_press <= 1'b0;
    end else begin
        debounce_cnt_prev <= (debounce_cnt >= DEBOUNCE_CNT);  // �������Ƿ��ȶ�����
        key_state <= (debounce_cnt >= DEBOUNCE_CNT);          // ��ǰ�ȶ�״̬����=���£�
        
        // ���ڡ�������δ�ȶ�����ǰ�����ȶ���ʱ�����1�����ڵ�key_press�����δ�����
        key_press <= (debounce_cnt >= DEBOUNCE_CNT) && (!debounce_cnt_prev);
    end
end

endmodule