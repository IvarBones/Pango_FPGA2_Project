`timescale 1ns/1ns
module defect_four_points_no_error_tb();

// -------------------------- �źŶ��� --------------------------
reg                     pixclk_in;       // ����ʱ��
reg                     rst_n;           // ��λ������Ч��
reg                     bin2_vs;         // ��ͬ���ź�
reg                     bin2_de;         // ������Ч�ź�
reg                     bin2_data;       // ��ֵ���������ݣ�1=覴ã�0=������
reg [7:0]               cnt;             // �����������ڿ���ʱ��

// ģ������ź�
wire [10:0]             defect_p1_x;     // ����1-X��x_min��
wire [10:0]             defect_p1_y;     // ����1-Y
wire [10:0]             defect_p2_x;     // ����2-X��x_max��
wire [10:0]             defect_p2_y;     // ����2-Y
wire [10:0]             defect_p3_x;     // ����3-X
wire [10:0]             defect_p3_y;     // ����3-Y��y_min��
wire [10:0]             defect_p4_x;     // ����4-X
wire [10:0]             defect_p4_y;     // ����4-Y��y_max��
wire                    defect_valid;    // 覴���Ч��־
wire                    point_vs;        // �ӳٳ�ͬ��
wire                    point_de;        // �ӳ�������Ч

// -------------------------- ��ʼ����ʱ������ --------------------------
initial begin
    pixclk_in    <= 1'd0;
    rst_n        <= 1'd0;
    bin2_vs      <= 1'd0;
    bin2_de      <= 1'd0;
    bin2_data    <= 1'd0;
    cnt          <= 8'd0;

    #20  // ��λ20ns���ͷ�
    rst_n <= 1'd1;
end

// 50MHz����ʱ�ӣ�����10ns������matrix_tb����һ��
always #10 pixclk_in = ~pixclk_in;

// -------------------------- ����������ʱ�� --------------------------
// ������ѭ��������0~19������������������Ч�ͳ�ͬ���ź�
always @(posedge pixclk_in or negedge rst_n) begin
    if (!rst_n)
        cnt <= 8'd0;
    else if (cnt >= 8'd19)  // ������19�����㣬����20*10ns=200ns
        cnt <= 8'd0;
    else
        cnt <= cnt + 1'b1;
end

// -------------------------- ���������ź� --------------------------
// 1. ��ͬ���ź�bin2_vs��ÿ֡��ʼʱ��cnt=0������1��ʱ������
always @(posedge pixclk_in or negedge rst_n) begin
    if (!rst_n)
        bin2_vs <= 1'd0;
    else
        bin2_vs <= (cnt == 8'd0) ? 1'd1 : 1'd0;  // ֡��ʼ���
end

// 2. ������Ч�ź�bin2_de��cnt=1~15�ڼ���Ч��ģ����Чͼ������
always @(posedge pixclk_in or negedge rst_n) begin
    if (!rst_n)
        bin2_de <= 1'd0;
    else if (cnt >= 8'd1 && cnt <= 8'd15)  // ��Ч���ݴ���
        bin2_de <= 1'd1;
    else
        bin2_de <= 1'd0;
end

// 3. ��ֵ��覴�����bin2_data��ģ��һ������覴�����
// 覴�λ�ã�����Ч���ݴ����ڣ�cnt=3~10���з������м���������3λ��=1~3���з���
reg [2:0] row_cnt;  // �м�������0~7ѭ����ģ��ͼ���У�
always @(posedge pixclk_in or negedge rst_n) begin
    if (!rst_n) begin
        row_cnt <= 3'd0;
        bin2_data <= 1'd0;
    end else begin
        // �м�������ÿ֡��20��ʱ�ӣ�ѭ��һ��
        row_cnt <= (cnt == 8'd19) ? row_cnt + 1'b1 : row_cnt;

        // 覴�������1~3����3~10��bin2_data=1��
        if (bin2_de) begin  // ��������Чʱ����覴�
            bin2_data <= (row_cnt >= 3'd1 && row_cnt <= 3'd3) 
                      && (cnt >= 8'd3 && cnt <= 8'd10) ? 1'd1 : 1'd0;
        end else begin
            bin2_data <= 1'd0;
        end
    end
end

// -------------------------- ʵ����������ģ�� --------------------------
// ������С�ߴ�ͼ��5x5�����ӿ�����ٶ�
defect_four_points_no_error#(
    .IMG_WIDTH    (11'd5),    // ͼ����5����0~4��
    .IMG_HEIGHT   (11'd5),    // ͼ��߶�5����0~4��
    .COORD_WID    (11),       // ����λ��11
    .DELAY_CYCLES (1)         // �ӳ�����1
) u_defect_four_points_no_error (
    .pixclk_in    (pixclk_in),
    .rstn_out     (rst_n),
    .bin2_vs      (bin2_vs),
    .bin2_de      (bin2_de),
    .bin2_data    (bin2_data),
    .defect_p1_x  (defect_p1_x),
    .defect_p1_y  (defect_p1_y),
    .defect_p2_x  (defect_p2_x),
    .defect_p2_y  (defect_p2_y),
    .defect_p3_x  (defect_p3_x),
    .defect_p3_y  (defect_p3_y),
    .defect_p4_x  (defect_p4_x),
    .defect_p4_y  (defect_p4_y),
    .defect_valid (defect_valid),
    .point_vs     (point_vs),
    .point_de     (point_de)
);

endmodule