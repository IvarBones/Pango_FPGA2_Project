module box_merger #(
    parameter MAX_BOX_NUM = 10,
    parameter BOX_WIDTH   = 38
)(
    input  wire clk,
    input  wire rst_n,

    input  wire vs_in,                 // ֡ͬ��
    input  wire eoc_in,                // box��Ч����
    input  wire [BOX_WIDTH-1:0] box_in,

    output reg  [3:0] box_count_out,   // ��Ч box �� (0~10)
    output wire [MAX_BOX_NUM*BOX_WIDTH-1:0] box_all_out
);

    // ==============================
    // 10 �������Ĵ���
    // ==============================
    reg [BOX_WIDTH-1:0] box0;
    reg [BOX_WIDTH-1:0] box1;
    reg [BOX_WIDTH-1:0] box2;
    reg [BOX_WIDTH-1:0] box3;
    reg [BOX_WIDTH-1:0] box4;
    reg [BOX_WIDTH-1:0] box5;
    reg [BOX_WIDTH-1:0] box6;
    reg [BOX_WIDTH-1:0] box7;
    reg [BOX_WIDTH-1:0] box8;
    reg [BOX_WIDTH-1:0] box9;

    reg [3:0] box_count; // 0~10

    // ==============================
    // д�� / �����߼�
    // ==============================
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            box_count <= 4'd0;
            // box0~box9 �����㣬����ͼ�����������/��ʧ����
        end
        else if(vs_in) begin
            // ��֡��ʼ��ֻ�������������ʷ����
            box_count <= 4'd0;
        end
        else if(eoc_in && box_count < MAX_BOX_NUM) begin
            case(box_count)
                4'd0: box0 <= box_in;
                4'd1: box1 <= box_in;
                4'd2: box2 <= box_in;
                4'd3: box3 <= box_in;
                4'd4: box4 <= box_in;
                4'd5: box5 <= box_in;
                4'd6: box6 <= box_in;
                4'd7: box7 <= box_in;
                4'd8: box8 <= box_in;
                4'd9: box9 <= box_in;
            endcase
            box_count <= box_count + 1'b1;
        end
    end

    // ��� box ����ͬ��������ɣ�
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n)
            box_count_out <= 4'd0;
        else if(vs_in)
            box_count_out <= box_count;
    end

    // ƴ�ӳɱ�ƽ�����˳��Ϊ box0 �����λ
    assign box_all_out = {
        box9, box8, box7, box6, box5,
        box4, box3, box2, box1, box0
    };

endmodule
