module binarization(
    input               clk             ,   
    input               rst_n           ,   

    input               vsync_in        ,   // ���볡ͬ��
    input               hsync_in        ,   // ������ͬ��
    input               de_in           ,   // ����������Ч
    input   [7:0]       y_in            ,   // ������������
    input   [7:0]       bin_threshold   ,   // ��������ֵ����̬��ֵ�����԰������ƣ�

    output              vsync_out       ,   // �����ͬ�����ӳ�1�ģ�
    output              hsync_out       ,   // �����ͬ�����ӳ�1�ģ�
    output              de_out          ,   // ���������Ч���ӳ�1�ģ�
    output   reg        pix                // ��ֵ�����
);

// �Ĵ������壨ͬ���ź��ã�
reg    vsync_in_d;
reg    hsync_in_d;
reg    de_in_d   ;

// ���ͬ���źţ����ֵ��������룬�ӳ�1�ģ�
assign  vsync_out = vsync_in_d  ;
assign  hsync_out = hsync_in_d  ;
assign  de_out    = de_in_d     ;

// ��ֵ���߼���ʹ�ö�̬��ֵ��
always @(posedge clk or negedge rst_n) begin
    if(!rst_n)
        pix <= 1'b0;
    else if(de_in)  // ����������Чʱ����
        pix <= (y_in > bin_threshold) ? 1'b1 : 1'b0;  // ��̬��ֵ�ж�
    else
        pix <= 1'b0;  // ��Ч�������0
end

// ͬ���ź��ӳ�1�ģ����ֵ�����ʱ����룩
always@(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        vsync_in_d <= 1'd0;
        hsync_in_d <= 1'd0;
        de_in_d    <= 1'd0;
    end
    else begin
        vsync_in_d <= vsync_in;
        hsync_in_d <= hsync_in;
        de_in_d    <= de_in   ;
    end
end

endmodule